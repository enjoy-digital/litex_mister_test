`define BUILD_DATE "20230412"
`define XILINX 1
`define MISTER_DEBUG_NOHDMI 1
`define MISTER_DOWNSCALE_NN 1
`define MISTER_DISABLE_YC 1
`define MISTER_DISABLE_ALSA 1
